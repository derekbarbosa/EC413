module Verification_64bit (sumv, a, b, c_in);

	input [63:0] a;
	input [63:0] b;
	input c_in;

	output [63:0]sumv; 

	assign {sumv} = a + b + c_in;

endmodule